module dataMEM_test();

reg clk, rst, E, RW; 
reg [63:0] A;
reg [63:0] B; 
output [31:0] O; 
reg [31:0] mem [0:65535];

dataMEM DUT(clk, rst, A, B, E, RW, O); 

initial
begin
    $display("Data Memory");
    $display(" ");
    $display("Test 1");
    clk <= 0;
    clk <= 1;

    rst <= 1;
    E <= 1;
    RW <= 0;
    A = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    B = 64'b0000000000000000000000000000000000011000000000110011111110000000;
    #100
    $display("Output = %b", O);


    $display(" ");
    $display("Test 2");
    clk <= 0;
    clk <= 1;

    rst <= 0;
    E <= 0;
    RW <= 0;
    A = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    B = 64'b0000000000000000000000011000000100000000000000111111111110000000;
    #100
    $display("Output = %b", O);


    $display(" ");
    $display("Test 3");
    clk <= 0;
    clk <= 1;
    
    rst <= 1;
    E <= 1;
    RW <= 0;
    A = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    B = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    #100
    $display("Output = %b", O);

end

endmodule
