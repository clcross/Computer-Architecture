// got help from sammy T
module registerfile (clk, rst, read1, read2, writeto, writedat, writeenable, out1, out2);
    input writeenable, clk, rst;
    input [4:0] read1; 
    input [4:0] read2; 
    input [4:0] writeto;
    input [63:0] writedat;
    output [63:0] out1, out2;

    reg [31:0] RF [63:0];

    assign #4 out1 = RF[read1];
    assign #4 out2 = RF[read2];

    always @(posedge clk)
    begin
        if (writeenable) RF[writeto] <= writedat;
            $display("regfile: %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[0], RF[1], RF[2], RF[3], RF[4], RF[5], RF[6], RF[7]);
            $display("         %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[8], RF[9], RF[10], RF[11], RF[12], RF[13], RF[14], RF[15]);
            $display("         %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[16], RF[17], RF[18], RF[19], RF[20], RF[21], RF[22], RF[23]);
            $display("         %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[24], RF[25], RF[26], RF[27], RF[28], RF[29], RF[30], RF[31]);
            $display("         %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[32], RF[33], RF[34], RF[35], RF[36], RF[37], RF[38], RF[39]);
            $display("         %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[40], RF[41], RF[42], RF[43], RF[44], RF[45], RF[46], RF[47]);
            $display("         %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[48], RF[49], RF[50], RF[51], RF[52], RF[53], RF[54], RF[55]);
            $display("         %h, %h, %h, %h, %h, %h, %h, %h,", 
                RF[56], RF[57], RF[58], RF[59], RF[60], RF[61], RF[62], RF[63]);
    end

    always @(posedge rst)
    begin
        RF[0] <= 64'h0000000000000000;
        RF[1] <= 64'h0000000000000000;
        RF[2] <= 64'h0000000000000000;
        RF[3] <= 64'h0000000000000000;
        RF[4] <= 64'h0000000000000000;
        RF[5] <= 64'h0000000000000000;
        RF[6] <= 64'h0000000000000000;
        RF[7] <= 64'h0000000000000000;
        RF[8] <= 64'h0000000000000000;
        RF[9] <= 64'h0000000000000000;
        RF[10] <= 64'h0000000000000000;
        RF[11] <= 64'h0000000000000000;
        RF[12] <= 64'h0000000000000000;
        RF[13] <= 64'h0000000000000000;
        RF[14] <= 64'h0000000000000000;
        RF[15] <= 64'h0000000000000000;
        RF[16] <= 64'h0000000000000000;
        RF[17] <= 64'h0000000000000000;
        RF[18] <= 64'h0000000000000000;
        RF[19] <= 64'h0000000000000000;
        RF[20] <= 64'h0000000000000000;
        RF[21] <= 64'h0000000000000000;
        RF[22] <= 64'h0000000000000000;
        RF[23] <= 64'h0000000000000000;
        RF[24] <= 64'h0000000000000000;
        RF[25] <= 64'h0000000000000000;
        RF[26] <= 64'h0000000000000000;
        RF[27] <= 64'h0000000000000000;
        RF[28] <= 64'h0000000000000000;
        RF[29] <= 64'h0000000000000000;
        RF[30] <= 64'h0000000000000000;
        RF[31] <= 64'h0000000000000000;
        RF[32] <= 64'h0000000000000000;
        RF[33] <= 64'h0000000000000000;
        RF[34] <= 64'h0000000000000000;
        RF[35] <= 64'h0000000000000000;
        RF[36] <= 64'h0000000000000000;
        RF[37] <= 64'h0000000000000000;
        RF[38] <= 64'h0000000000000000;
        RF[39] <= 64'h0000000000000000;
        RF[40] <= 64'h0000000000000000;
        RF[41] <= 64'h0000000000000000;
        RF[42] <= 64'h0000000000000000;
        RF[43] <= 64'h0000000000000000;
        RF[44] <= 64'h0000000000000000;
        RF[45] <= 64'h0000000000000000;
        RF[46] <= 64'h0000000000000000;
        RF[47] <= 64'h0000000000000000;
        RF[48] <= 64'h0000000000000000;
        RF[49] <= 64'h0000000000000000;
        RF[50] <= 64'h0000000000000000;
        RF[51] <= 64'h0000000000000000;
        RF[52] <= 64'h0000000000000000;
        RF[53] <= 64'h0000000000000000;
        RF[54] <= 64'h0000000000000000;
        RF[55] <= 64'h0000000000000000;
        RF[56] <= 64'h0000000000000000;
        RF[57] <= 64'h0000000000000000;
        RF[58] <= 64'h0000000000000000;
        RF[59] <= 64'h0000000000000000;
        RF[60] <= 64'h0000000000000000;
        RF[61] <= 64'h0000000000000000;
        RF[62] <= 64'h0000000000000000;
        RF[63] <= 64'h0000000000000000;
    end
endmodule

// module registerfile (clk, rst, read1, read2, writeto, writedat, writeenable, out1, out2); 
//     input writeenable, clk, rst; 
//     input [4:0] read1; 
//     input [4:0] read2; 
//     input [4:0] writeto; 
//     input [63:0] writedat; 
//     output [63:0] out1, out2; 
//     // 32 bit registers x 32 
//     reg [63:0] RF [31:0];

//     assign #2 out1 = RF[read1];
//     assign #2 out2 = RF[read2];

//     always @ (negedge clk) 
//     begin
//         if(writeenable)
//         if (writeto != 4'd31)
//             RF[writeto] <= #3 writedat;
//         else 
//             RF[0] <= #3 'd0; 
//     end

// endmodule